../../../src/04-sequential-logic/sum_reduce/sum_reduce.sv