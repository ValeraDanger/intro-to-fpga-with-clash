../../../src/01-intro-to-simulation/hello_world.sv