module hello_world;
  initial begin
    $display("Hello world!");
    $finish;
  end
endmodule
