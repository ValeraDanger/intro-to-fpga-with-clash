../../../src/02-combination-logic/testbenches/adder_1_bit_tb.sv