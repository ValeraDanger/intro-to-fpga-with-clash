../../../src/03-principles-of-constructor/adder_multibits_bitvectors.sv