../../../src/02-adder/adder_plus_1_bit.sv