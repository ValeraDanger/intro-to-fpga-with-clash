../../../src/02-combination-logic/adder_plus_1_bit.sv