module adder_multibits_int(
  input int a,
  input int b,
  output int sum
);
  assign sum = a + b;
endmodule
