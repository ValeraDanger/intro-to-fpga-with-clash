../../../src/02-adder/testbenches/adder_1_bit_tb.sv