../../../src/02-combination-logic/adder_logic_1_bit_tb.sv