../../../src/02-adder/adder_logic_1_bit.sv