../../../src/03-principles-of-constructor/adder_reuse_without_generate.sv