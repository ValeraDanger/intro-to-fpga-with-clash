../../../src/01-basic-environment/hello_world.sv